
`ifndef _UART_DEFINES_
`define _UART_DEFINES_


`define STOP_BITS_ONE            1
`define STOP_BITS_ONE_POINT_FIVE 2
`define STOP_BITS_TWO            3 

`define PARITY_NONE 1
`define PARITY_ODD  2
`define PARITY_EVEN 3          


`endif